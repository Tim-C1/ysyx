module ifu (
    input pc,
    output [63:0] inst
)

// pass
